blueBox.png ballBlue
yellowBall.png ballYellow
blueBoxCrouch.png ballCrouch
redBox.png box
redSlab.png slab
ground.png ground
bullet.png bullet
wall.png wall
heal.png healCollect
hpUp.png hpUpCollect
dmgUp.png dmgUpCollect
fasterShots.png fasterShotsCollect
fasterShooting.png fasterShootingCollect
noReload.png noReloadCollect
health.png healthBar