Player{
    ObjectProperties{
        position 89 -1
        name player2
        texture humanMale
    }
    PhysicObjectProperties{
        type dynamic
        shape circle
        friction 0.1
        density 1
    }
    EntityProperties{
        maxHP 10
        HP 10
        jumpHeight 300
        movementSpeed 10
        EQ{
            rodBrown 10 0
            bow 1 0
        }
    }
    PlayerProperties{
        textureBase humanMale
        textureHair aragornHair
        textureBoots bootsMiddleGray
        textureLegs legArmor0
        textureGloves gloveBrown
        textureBody aragornBody
        textureCloak cloackBlack
    }
}