Player{
    ObjectProperties{
        position 89 -1
        name player2
        texture humanMale
    }
    PhysicObjectProperties{
        type dynamic
        shape circle
        friction 0.1
        density 1
    }
    EntityProperties{
        maxHP 250
        HP 250
        jumpHeight 300
        movementSpeed 10
        equiped 1
        EQ{
            rodBrown 10 0
            bow 1 0
            laserRod 50 0
        }
    }
    PlayerProperties{
        textureBase humanMale
        textureHair aragornHair
        textureBoots bootsMiddleGray
        textureLegs legArmor0
        textureGloves gloveBrown
        textureBody aragornBody
        textureCloak cloackBlack
    }
}
