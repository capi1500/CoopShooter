Player{
	ObjectProperties{
		position 89 -0.974279
		name player2
		texture humanMale
	}
	PhysicObjectProperties{
		type dynamic
		shape circle
		density 1
		friction 0.1
		angle 0
		velocity 0 0
	}
	EntityProperties{
		maxHP 250
		HP 250
		jumpHeight 300
		movementSpeed 10
		isFacingLeft true
		equiped 1
		EQ{
			rodBrown 10 7346
			bow 1 7346
			laserRod 50 7346
			nothing 0
			nothing 0
		}
	}
	PlayerProperties{
		textureBase humanMale
		textureHair aragornHair
		textureBoots bootsMiddleGray
		textureLegs legArmor0
		textureGloves gloveBrown
		textureBody aragornBody
		textureHandRight bowEquiped
		textureCloak cloackBlack
		textureBeard nothing
	}
}
