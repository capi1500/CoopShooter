Player{
	ObjectProperties{
		position 8.72241 -2.97479
		name player1
		texture humanMale
	}
	PhysicObjectProperties{
		type dynamic
		shape circle
		density 1
		friction 0.1
		angle 0
		velocity -14.9815 0
	}
	EntityProperties{
		maxHP 250
		HP 250
		jumpHeight 300
		movementSpeed 10
		isFacingLeft false
		equiped 1
		EQ{
			dagger 1 7346
			laserRod 50 368
			nothing 0
			nothing 0
			nothing 0
		}
	}
	PlayerProperties{
		textureBase humanMale
		textureHair longWhiteHair
		textureBoots bootsMiddleGray
		textureLegs nothing
		textureGloves nothing
		textureBody gandalfBody
		textureHandRight laserRodEquiped
		textureCloak cloackGray
		textureBeard nothing
	}
}
