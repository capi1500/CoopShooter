blockSize 32 32
startPos 0 0
Temp ground {
    ObjectProperties{
        position -1 0
    }
}
Temp ground {
    ObjectProperties{
        position 0 0
    }
}
Temp ground {
    ObjectProperties{
        position 1 0
    }
}
Temp ground {
    ObjectProperties{
        position 2 0
    }
}
Temp ground {
    ObjectProperties{
        position 3 0
    }
}
Temp ground {
    ObjectProperties{
        position 4 0
    }
}
Temp ground {
    ObjectProperties{
        position 5 0
    }
}
Temp ground {
    ObjectProperties{
        position 6 0
    }
}
Temp ground {
    ObjectProperties{
        position 7 0
    }
}
Temp ground {
    ObjectProperties{
        position 8 0
    }
}
Temp ground {
    ObjectProperties{
        position 9 0
    }
}
Temp ground {
    ObjectProperties{
        position 10 0
    }
}
Temp ground {
    ObjectProperties{
        position 11 0
    }
}
Temp ground {
    ObjectProperties{
        position 12 0
    }
}
Temp ground {
    ObjectProperties{
        position 13 0
    }
}
Temp ground {
    ObjectProperties{
        position 14 0
    }
}
Temp ground {
    ObjectProperties{
        position 15 0
    }
}
Temp ground {
    ObjectProperties{
        position 16 0
    }
}
Temp ground {
    ObjectProperties{
        position 17 0
    }
}
Temp ground {
    ObjectProperties{
        position 18 0
    }
}
Temp ground {
    ObjectProperties{
        position 19 0
    }
}
Temp ground {
    ObjectProperties{
        position 20 0
    }
}
Temp ground {
    ObjectProperties{
        position 21 0
    }
}
Temp ground {
    ObjectProperties{
        position 22 0
    }
}
Temp ground {
    ObjectProperties{
        position 23 0
    }
}
Temp ground {
    ObjectProperties{
        position 24 0
    }
}
Temp ground {
    ObjectProperties{
        position 25 0
    }
}
Temp ground {
    ObjectProperties{
        position 26 0
    }
}
Temp ground {
    ObjectProperties{
        position 27 0
    }
}
Temp ground {
    ObjectProperties{
        position 28 0
    }
}
Temp ground {
    ObjectProperties{
        position 29 0
    }
}
Temp ground {
    ObjectProperties{
        position -1 -1
    }
}
Temp ground {
    ObjectProperties{
        position -1 -2
    }
}
Temp ground {
    ObjectProperties{
        position -1 -3
    }
}
Temp ground {
    ObjectProperties{
        position -1 -4
    }
}
Temp ground {
    ObjectProperties{
        position -1 -5
    }
}
Temp ground {
    ObjectProperties{
        position -1 -6
    }
}
Temp ground {
    ObjectProperties{
        position -1 -7
    }
}
Temp ground {
    ObjectProperties{
        position -1 -8
    }
}
Temp ground {
    ObjectProperties{
        position -1 -9
    }
}
Temp ground {
    ObjectProperties{
        position -1 -10
    }
}
Temp groundSlab {
    ObjectProperties{
        position 2 -1.75
    }
}
Temp ground {
    ObjectProperties{
        position 2 -1
    }
}
Temp groundSlab {
    ObjectProperties{
        position 0 -3.75
    }
}
Temp groundSlab {
    ObjectProperties{
        position 1 -3.75
    }
}
Temp groundSlab {
    ObjectProperties{
        position 2 -3.75
    }
}
Temp groundSlab {
    ObjectProperties{
        position 3 -1.75
    }
}
Temp groundSlab {
    ObjectProperties{
        position 5 -3
    }
}
Temp groundSlab {
    ObjectProperties{
        position  6 -3
    }
}
Temp groundSlab {
    ObjectProperties{
        position 7 -3
    }
}
Temp groundSlab {
    ObjectProperties{
        position 8 -5
    }
}
Temp groundSlab {
    ObjectProperties{
        position 9 -5
    }
}
Temp ground {
    ObjectProperties{
        position 9 -2
    }
}
Temp ground {
    ObjectProperties{
        position 6 -1
    }
}
Temp groundSlab {
    ObjectProperties{
        position 11.5 -4.25
    }
}
Temp groundSlab {
    ObjectProperties{
        position 12.5 -4.25
    }
}
Temp groundSlab {
    ObjectProperties{
        position 10 -2.25
    }
}
Temp groundSlab {
    ObjectProperties{
        position 12 -0.75
    }
}
Temp ground {
    ObjectProperties{
        position 13 -2.5
    }
}
Temp ground {
    ObjectProperties{
        position 14.5 -6
    }
}
Temp ground {
    ObjectProperties{
        position 14.5 -7
    }
}
Temp groundSlab {
    ObjectProperties{
        position 13 -0.75
    }
}
Temp groundSlab {
    ObjectProperties{
        position 14 -0.75
    }
}
Temp groundSlab {
    ObjectProperties{
        position 15 -0.75
    }
}
Temp groundSlab {
    ObjectProperties{
        position 16 -0.75
    }
}
Temp ground {
    ObjectProperties{
        position 16 -2.5
    }
}
Temp groundSlab {
    ObjectProperties{
        position 17 -0.75
    }
}
Temp groundSlab {
    ObjectProperties{
        position 17 -0.75
    }
}
Temp groundSlab {
    ObjectProperties{
        position 19 -2.25
    }
}
Temp groundSlab {
    ObjectProperties{
        position 16.5 -4.25
    }
}
Temp groundSlab {
    ObjectProperties{
        position 17.5 -4.25
    }
}
Temp groundSlab {
    ObjectProperties{
        position 27 -1.75
    }
}
Temp ground {
    ObjectProperties{
        position 27 -1
    }
}
Temp groundSlab {
    ObjectProperties{
        position 29 -3.75
    }
}
Temp groundSlab {
    ObjectProperties{
        position 28 -3.75
    }
}
Temp groundSlab {
    ObjectProperties{
        position 27 -3.75
    }
}
Temp groundSlab {
    ObjectProperties{
        position 26 -1.75
    }
}
Temp groundSlab {
    ObjectProperties{
        position 24 -3
    }
}
Temp groundSlab {
    ObjectProperties{
        position 23 -3
    }
}
Temp groundSlab {
    ObjectProperties{
        position 22 -3
    }
}
Temp groundSlab {
    ObjectProperties{
        position 21 -5
    }
}
Temp groundSlab {
    ObjectProperties{
        position 20 -5
    }
}
Temp ground {
    ObjectProperties{
        position 20 -2
    }
}
Temp ground {
    ObjectProperties{
        position 23 -1
    }
}
Spawn{
    position 2 -2.5
}
Spawn{
    position 27 -2.5
}
Spawn{
    position 10 -3
}
Spawn{
    position 19 -3
}