Weapon{
	ObjectProperties{
		position -0.969697 -0.969697
		name bow
		texture bow
	}
	ItemProperties{
		amount -950389584
		isWorldObject true
		textureOnEquip bowEquiped
	}
	WeaponProperties{
		attackDelay 500
		bulletSpeed 1000
		dmg 6
		reloadSpeed 500
		maxAmmo 1
		ammo 1
		bulletTexture arrow
		bulletDistance 50
		reloading false
	}
}
Item{
	ObjectProperties{
		position 0 0
		name nothing
		texture }
	}
	ItemProperties{
		amount 1
		isWorldObject false
		textureOnEquip nothing
	}
}
Weapon{
	ObjectProperties{
		position -0.969697 -0.969697
		name rodBrown
		texture rodBrown
	}
	ItemProperties{
		amount -950495088
		isWorldObject true
		textureOnEquip rodBrownEquiped
	}
	WeaponProperties{
		attackDelay 350
		bulletSpeed 1000
		dmg 2
		reloadSpeed 3000
		maxAmmo 10
		ammo 10
		bulletTexture laser
		bulletDistance 20
		reloading false
	}
}
Weapon{
	ObjectProperties{
		position -0.969697 -0.969697
		name staff
		texture staff
	}
	ItemProperties{
		amount -950495184
		isWorldObject true
		textureOnEquip staffRubyEquiped
	}
	WeaponProperties{
		attackDelay 300
		bulletSpeed 1000
		dmg 2
		reloadSpeed 3000
		maxAmmo 20
		ammo 20
		bulletTexture fireball
		bulletDistance 30
		reloading false
	}
}
