Weapon{
    ObjectProperties{
        name bow
        texture bow
    }
    ItemProperties{
        ammount 1
        worldObject false
    }
    WeaponProperties{
        attackDelay 250
        bulletSpeed 50
        dmg 2
        reloadSpeed 3000
        maxAmmo 15
        bulletTexture arrow
        bulletDistance 50
    }
}
Weapon{
    ObjectProperties{
        name laserPistol
        texture laserPistol
    }
    ItemProperties{
        ammount 1
        worldObject false
    }
    WeaponProperties{
        attackDelay 350
        bulletSpeed 50
        dmg 4
        reloadSpeed 2000
        maxAmmo 10
        bulletTexture laser
        bulletDistance 20
    }
}
Weapon{
    ObjectProperties{
        name staff
        texture staff
    }
    ItemProperties{
        ammount 1
        worldObject false
    }
    WeaponProperties{
        attackDelay 300
        bulletSpeed 50
        dmg 2
        reloadSpeed 3000
        maxAmmo 20
        bulletTexture fireball
        bulletDistance 30
    }
}