Weapon{
    ObjectProperties{
        name bow
        texture bow
    }
    ItemProperties{
        ammount 1
        worldObject false
        textureOnEquip bowEquiped
    }
    WeaponProperties{
        attackDelay 600
        bulletSpeed 1000
        dmg 7
        reloadSpeed 1000
        maxAmmo 1
        bulletTexture arrow
        bulletDistance 55
        shotSound arrow
    }
}
Weapon{
    ObjectProperties{
        name rodBrown
        texture rodBrown
    }
    ItemProperties{
        ammount 1
        worldObject false
        textureOnEquip rodBrownEquiped
    }
    WeaponProperties{
        attackDelay 250
        bulletSpeed 1000
        dmg 2
        reloadSpeed 1000
        maxAmmo 10
        bulletTexture laser
        bulletDistance 10
        shotSound magicMissle
    }
}
Weapon{
    ObjectProperties{
        name staff
        texture staff
    }
    ItemProperties{
        ammount 1
        worldObject false
        textureOnEquip staffRubyEquiped
    }
    WeaponProperties{
        attackDelay 400
        bulletSpeed 1000
        dmg 3
        reloadSpeed 3000
        maxAmmo 20
        bulletTexture fireball
        bulletDistance 25
        shotSound fireball
    }
}
Weapon{
    ObjectProperties{
        name dagger
        texture dagger
    }
    ItemProperties{
        ammount 1
        worldObject false
        textureOnEquip daggerEquiped
    }
    WeaponProperties{
        attackDelay 1000
        bulletSpeed 500
        dmg 100
        reloadSpeed 1000
        maxAmmo 1
        bulletTexture transparent
        bulletDistance 0.01
        shotSound arrow
    }
}
Weapon{
    ObjectProperties{
        name laserRod
        texture laserRod
    }
    ItemProperties{
        ammount 1
        worldObject false
        textureOnEquip laserRodEquiped
    }
    WeaponProperties{
        attackDelay 25
        bulletSpeed 350
        dmg 1
        reloadSpeed 3000
        maxAmmo 50
        bulletTexture laserBall
        bulletDistance 2
        shotSound laserBall
    }
}
Item{
    ObjectProperties{
        name nothing
    }
    ItemProperties{
        ammount 0
        worldObject false
    }
}
