Player{
	ObjectProperties{
		position 54.7403 -3.65942
		name player2
		texture humanMale
	}
	PhysicObjectProperties{
		type dynamic
		shape circle
		density 1
		friction 0.1
		angle 0
		velocity -59.429 -42.9434
	}
	EntityProperties{
		maxHP 10
		HP 0
		jumpHeight 300
		movementSpeed 10
		isFacingLeft false
		equiped 2
		EQ{
			rodBrown 1 10765
			bow 1 4003
			rodBrown 7 5660
			nothing 0
			nothing 0
		}
	}
	PlayerProperties{
		textureBase humanMale
		textureHair aragornHair
		textureBoots bootsMiddleGray
		textureLegs legArmor0
		textureGloves gloveBrown
		textureBody aragornBody
		textureHandRight rodBrownEquiped
		textureCloak cloackBlack
		textureBeard nothing
	}
}
