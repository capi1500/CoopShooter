Assets/Textures/ammo.png ammoBar 0 0 28 64 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/player/body/aragorn.png aragornBody 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/player/hair/aragorn.png aragornHair 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/effect/arrow_2.png arrow 5 13 22 6 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/player/boots/middle_gray.png bootsMiddleGray 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/item/weapon/ranged/longbow_1.png bow 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/player/hand_right/bow.png bowEquiped 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/dungeon/wall/stone_brick_1.png box 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/player/cloak/black.png cloackBlack 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/player/cloak/gray.png cloackGray 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/item/potion/golden.png dmgUp 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/misc/slot.png eqItem 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/misc/slot_vehumet.png eqItemSelected 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/item/potion/ruby_new.png fasterShooting 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/item/potion/brilliant_blue_new.png fasterShots 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/effect/flame_0.png fireball 9 9 14 14 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/player/body/gandalf_g.png gandalfBody 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/player/gloves/glove_brown.png gloveBrown 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/item/potion/magenta_new.png heal 0 0 32 32 ;
Assets/Textures/health.png healthBar 0 0 28 64 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/item/potion/bubbly.png hpUp 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/player/base/human_male.png humanMale 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/effect/icicle_2.png laser 2 13 28 6 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/player/legs/leg_armor_0.png legArmor0 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/player/beard/long_white.png longWhiteBeard 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/player/hair/long_white.png longWhiteHair 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/item/potion/white_new.png noReload 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/item/rod/rod_1_new.png rodBrown 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/player/hand_right/rod_brown_new.png rodBrownEquiped 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/dungeon/wall/stone_brick_1.png slab 0 0 32 16 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/item/wand/gem_gold_new.png staff 0 0 32 32 ;
Assets/Textures/Dungeon_Crawl_Stone_Soup/player/hand_right/staff_ruby.png staffRubyEquiped 0 0 32 32 ;
Assets/Textures/blackScr.png blackScr ;
Assets/Textures/blackScr2.png blackScr2 ;
Assets/Textures/test.png logo ;
