Weapon{
    ObjectProperties{
        name bow
        texture bow
    }
    ItemProperties{
        ammount 1
        worldObject false
        textureOnEquip bowEquiped
        spawnable true
    }
    WeaponProperties{
        attackDelay 600
        bulletSpeed 1000
        dmg 70
        reloadSpeed 1000
        maxAmmo 1
        bulletTexture arrow
        bulletDistance 55
        shotSound arrow
    }
}
Weapon{
    ObjectProperties{
        name rodBrown
        texture rodBrown
    }
    ItemProperties{
        ammount 1
        worldObject false
        textureOnEquip rodBrownEquiped
        spawnable true
    }
    WeaponProperties{
        attackDelay 250
        bulletSpeed 1000
        dmg 20
        reloadSpeed 1000
        maxAmmo 10
        bulletTexture laser
        bulletDistance 10
        shotSound magicMissle
    }
}
Weapon{
    ObjectProperties{
        name staff
        texture staff
    }
    ItemProperties{
        ammount 1
        worldObject false
        textureOnEquip staffRubyEquiped
        spawnable true
    }
    WeaponProperties{
        attackDelay 400
        bulletSpeed 1000
        dmg 30
        reloadSpeed 3000
        maxAmmo 20
        bulletTexture fireball
        bulletDistance 25
        shotSound fireball
    }
}
Weapon{
    ObjectProperties{
        name dagger
        texture dagger
    }
    ItemProperties{
        ammount 1
        worldObject false
        textureOnEquip daggerEquiped
        spawnable true
    }
    WeaponProperties{
        attackDelay 1000
        bulletSpeed 500
        dmg 125
        reloadSpeed 1000
        maxAmmo 1
        bulletTexture transparent
        bulletDistance 0.01
        shotSound arrow
    }
}
Weapon{
    ObjectProperties{
        name ohBabeItsTripleDagger
        texture ohBabeItsTripleDagger
    }
    ItemProperties{
        ammount 1
        worldObject false
        textureOnEquip ohBabeItsTripleDaggerEquiped
        spawnable true
    }
    WeaponProperties{
        attackDelay 1000
        bulletSpeed 500
        dmg 1000
        reloadSpeed 1000
        maxAmmo 1
        bulletTexture transparent
        bulletDistance 0.01
        shotSound arrow
    }
}
Weapon{
    ObjectProperties{
        name laserRod
        texture laserRod
    }
    ItemProperties{
        ammount 1
        worldObject false
        textureOnEquip laserRodEquiped
        spawnable true
    }
    WeaponProperties{
        attackDelay 25
        bulletSpeed 350
        dmg 5
        reloadSpeed 3000
        maxAmmo 50
        bulletTexture laserBall
        bulletDistance 2
        shotSound laserBall
    }
}
Item{
    ObjectProperties{
        name nothing
    }
    ItemProperties{
        ammount 0
        worldObject false
    }
}