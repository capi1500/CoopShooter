Weapon{
	ObjectProperties{
		position -1.45455 -1.45455
		name bow
		texture bow
	}
	ItemProperties{
		amount 471676512
		isWorldObject true
		textureOnEquip bowEquiped
	}
	WeaponProperties{
		attackDelay 500
		bulletSpeed 1000
		dmg 6
		reloadSpeed 500
		maxAmmo 1
		ammo 1
		bulletTexture arrow
		bulletDistance 50
		reloading false
	}
}
Item{
	ObjectProperties{
		position 0 0
		name nothing
		texture }
	}
	ItemProperties{
		amount 1
		isWorldObject false
		textureOnEquip nothing
	}
}
Weapon{
	ObjectProperties{
		position -1.45455 -1.45455
		name rodBrown
		texture rodBrown
	}
	ItemProperties{
		amount 471571792
		isWorldObject true
		textureOnEquip rodBrownEquiped
	}
	WeaponProperties{
		attackDelay 350
		bulletSpeed 1000
		dmg 2
		reloadSpeed 3000
		maxAmmo 10
		ammo 10
		bulletTexture laser
		bulletDistance 20
		reloading false
	}
}
Weapon{
	ObjectProperties{
		position -1.45455 -1.45455
		name staff
		texture staff
	}
	ItemProperties{
		amount 471571696
		isWorldObject true
		textureOnEquip staffRubyEquiped
	}
	WeaponProperties{
		attackDelay 300
		bulletSpeed 1000
		dmg 2
		reloadSpeed 3000
		maxAmmo 20
		ammo 20
		bulletTexture fireball
		bulletDistance 30
		reloading false
	}
}
