arrow Assets/Audio/RPG-SFX/wood_02.ogg
collect Assets/Audio/BonusCube.ogg
eqChange Assets/Audio/RPG-SFX/misc_01.ogg
fireball Assets/Audio/RPG-SFX/spell_02.ogg
jump Assets/Audio/jump.ogg
magicMissle Assets/Audio/RPG-SFX/spell_01.ogg
menu Assets/Audio/menu.wav
