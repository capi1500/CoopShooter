Assets/Audio/RPG-SFX/wood_02.ogg arrow
Assets/Audio/BonusCube.ogg collect
Assets/Audio/RPG-SFX/misc_01.ogg eqChange
Assets/Audio/RPG-SFX/spell_02.ogg fireball
Assets/Audio/jump.ogg jump
Assets/Audio/RPG-SFX/spell_01.ogg magicMissle
Assets/Audio/menu.wav menu
