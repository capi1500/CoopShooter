wall.png box
slab.png slab
ground.png ground
wall.png wall
heal.png heal
hpUp.png hpUp
dmgUp.png dmgUp
fasterShots.png fasterShots
fasterShooting.png fasterShooting
noReload.png noReload
health.png healthBar
ammo.png ammoBar
battlemage.png mage
archer.png archer
arrow.png arrow
fireball.png fireball
bow.png bow
laserPistol.png laserPistol
sceptre.png staff
eqItem.png eqItem
eqItemSelected.png eqItemSelected
laser.png laser