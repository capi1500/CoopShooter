Player{
    ObjectProperties{
        position 1180 -35
        name player2
        texture archer
    }
    PhysicObjectProperties{
        type dynamic
        shape circle
        friction 0.1
        density 1
    }
    EntityProperties{
        maxHP 10
        HP 10
        jumpHeight 300
        movementSpeed 10
        EQ{
            assultRifle 1
        }
    }
}