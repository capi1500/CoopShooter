Player{
    ObjectProperties{
        position 89 -1
        name player2
        texture archer
    }
    PhysicObjectProperties{
        type dynamic
        shape circle
        friction 0.1
        density 1
    }
    EntityProperties{
        maxHP 10
        HP 10
        jumpHeight 300
        movementSpeed 10
        EQ{
            laserPistol 1
            bow 1
        }
    }
}