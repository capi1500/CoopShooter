Template{
    name ground
    WorldObject{
	    ObjectProperties{
	        texture box
	    }
	    PhysicObjectProperties{
            shape box
	    }
    }
}
Template{
    name groundSlab
    WorldObject{
	    ObjectProperties{
	        texture slab
	    }
	    PhysicObjectProperties{
            shape box
	    }
    }
}