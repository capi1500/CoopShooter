wall.gif box
slab.gif slab
ground.png ground
bullet.png bullet
wall.png wall
heal.png healCollect
hpUp.png hpUpCollect
dmgUp.png dmgUpCollect
fasterShots.png fasterShotsCollect
fasterShooting.png fasterShootingCollect
noReload.png noReloadCollect
health.png healthBar
ammo.png ammoBar
battlemage.gif mage
archer.gif archer
arrow.png arrow
fireball.gif fireball