blockSize 33 33
startPos 0 0
time 0.016523
Collectible{
	ObjectProperties{
		position 40 -3
		name collectible1320.000000--99.000000
		texture hpUp
	}
	PhysicObjectProperties{
		type kinematic
		shape circle
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	CollectibleProperties{
		what hpUp
		boostTime 0
	}
}
WorldObject{
	ObjectProperties{
		position -1 0
		name ground0
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 0 0
		name ground1
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 9 0
		name ground10
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 44 0
		name ground100
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 45 0
		name ground101
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 46 0
		name ground102
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 47 0
		name ground103
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 48 0
		name ground104
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 49 0
		name ground105
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 50 0
		name ground106
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 51 0
		name ground107
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 52 0
		name ground108
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 53 0
		name ground109
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 10 0
		name ground11
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 54 0
		name ground110
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 55 0
		name ground111
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 56 0
		name ground112
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 57 0
		name ground113
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 58 0
		name ground114
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 59 0
		name ground115
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 32 -1
		name ground117
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 11 0
		name ground12
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 39 -2
		name ground127
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 36 -1
		name ground128
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 12 0
		name ground13
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 43 -2.5
		name ground133
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 44.5 -6
		name ground134
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 44.5 -7
		name ground135
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 13 0
		name ground14
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 46 -2.5
		name ground140
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 57 -1
		name ground147
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 14 0
		name ground15
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 50 -2
		name ground157
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 53 -1
		name ground158
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 60 0
		name ground159
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 15 0
		name ground16
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 61 0
		name ground160
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 62 0
		name ground161
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 63 0
		name ground162
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 64 0
		name ground163
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 65 0
		name ground164
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 66 0
		name ground165
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 67 0
		name ground166
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 68 0
		name ground167
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 69 0
		name ground168
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 70 0
		name ground169
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 16 0
		name ground17
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 71 0
		name ground170
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 72 0
		name ground171
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 73 0
		name ground172
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 74 0
		name ground173
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 75 0
		name ground174
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 76 0
		name ground175
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 77 0
		name ground176
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 78 0
		name ground177
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 79 0
		name ground178
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 80 0
		name ground179
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 17 0
		name ground18
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 81 0
		name ground180
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 82 0
		name ground181
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 83 0
		name ground182
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 84 0
		name ground183
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 85 0
		name ground184
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 86 0
		name ground185
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 87 0
		name ground186
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 88 0
		name ground187
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 89 0
		name ground188
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 90 0
		name ground189
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 18 0
		name ground19
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 90 -1
		name ground190
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 90 -2
		name ground191
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 90 -3
		name ground192
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 90 -4
		name ground193
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 90 -5
		name ground194
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 90 -6
		name ground195
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 90 -7
		name ground196
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 90 -8
		name ground197
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 90 -9
		name ground198
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 90 -10
		name ground199
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 1 0
		name ground2
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 19 0
		name ground20
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 90 -11
		name ground200
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 62 -1
		name ground202
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 20 0
		name ground21
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 69 -2
		name ground212
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 66 -1
		name ground213
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 73 -2.5
		name ground218
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 74.5 -6
		name ground219
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 21 0
		name ground22
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 74.5 -7
		name ground220
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 76 -2.5
		name ground225
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 22 0
		name ground23
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 87 -1
		name ground232
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 23 0
		name ground24
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 80 -2
		name ground242
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 83 -1
		name ground243
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 24 0
		name ground25
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 25 0
		name ground26
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 26 0
		name ground27
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 27 0
		name ground28
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 28 0
		name ground29
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 2 0
		name ground3
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 29 0
		name ground30
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position -1 -1
		name ground31
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position -1 -2
		name ground32
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position -1 -3
		name ground33
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position -1 -4
		name ground34
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position -1 -5
		name ground35
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position -1 -6
		name ground36
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position -1 -7
		name ground37
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position -1 -8
		name ground38
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position -1 -9
		name ground39
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 3 0
		name ground4
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position -1 -10
		name ground40
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position -1 -11
		name ground41
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 2 -1
		name ground43
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 4 0
		name ground5
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 9 -2
		name ground53
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 6 -1
		name ground54
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 13 -2.5
		name ground59
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 5 0
		name ground6
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 14.5 -6
		name ground60
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 14.5 -7
		name ground61
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 16 -2.5
		name ground66
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 6 0
		name ground7
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 27 -1
		name ground73
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 7 0
		name ground8
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 20 -2
		name ground83
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 23 -1
		name ground84
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 29 0
		name ground85
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 30 0
		name ground86
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 31 0
		name ground87
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 32 0
		name ground88
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 33 0
		name ground89
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 8 0
		name ground9
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 34 0
		name ground90
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 35 0
		name ground91
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 36 0
		name ground92
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 37 0
		name ground93
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 38 0
		name ground94
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 39 0
		name ground95
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 40 0
		name ground96
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 41 0
		name ground97
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 42 0
		name ground98
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 43 0
		name ground99
		texture box
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 32 -1.75
		name groundSlab116
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 30 -3.75
		name groundSlab118
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 31 -3.75
		name groundSlab119
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 32 -3.75
		name groundSlab120
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 33 -1.75
		name groundSlab121
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 35 -3
		name groundSlab122
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 36 -3
		name groundSlab123
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 37 -3
		name groundSlab124
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 38 -5
		name groundSlab125
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 39 -5
		name groundSlab126
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 41.5 -4.25
		name groundSlab129
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 42.5 -4.25
		name groundSlab130
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 40 -2.25
		name groundSlab131
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 42 -0.75
		name groundSlab132
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 43 -0.75
		name groundSlab136
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 44 -0.75
		name groundSlab137
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 45 -0.75
		name groundSlab138
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 46 -0.75
		name groundSlab139
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 47 -0.75
		name groundSlab141
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 47 -0.75
		name groundSlab142
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 49 -2.25
		name groundSlab143
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 46.5 -4.25
		name groundSlab144
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 47.5 -4.25
		name groundSlab145
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 57 -1.75
		name groundSlab146
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 59 -3.75
		name groundSlab148
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 58 -3.75
		name groundSlab149
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 57 -3.75
		name groundSlab150
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 56 -1.75
		name groundSlab151
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 54 -3
		name groundSlab152
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 53 -3
		name groundSlab153
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 52 -3
		name groundSlab154
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 51 -5
		name groundSlab155
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 50 -5
		name groundSlab156
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 62 -1.75
		name groundSlab201
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 60 -3.75
		name groundSlab203
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 61 -3.75
		name groundSlab204
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 62 -3.75
		name groundSlab205
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 63 -1.75
		name groundSlab206
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 65 -3
		name groundSlab207
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 66 -3
		name groundSlab208
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 67 -3
		name groundSlab209
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 68 -5
		name groundSlab210
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 69 -5
		name groundSlab211
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 71.5 -4.25
		name groundSlab214
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 72.5 -4.25
		name groundSlab215
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 70 -2.25
		name groundSlab216
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 72 -0.75
		name groundSlab217
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 73 -0.75
		name groundSlab221
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 74 -0.75
		name groundSlab222
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 75 -0.75
		name groundSlab223
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 76 -0.75
		name groundSlab224
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 77 -0.75
		name groundSlab226
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 77 -0.75
		name groundSlab227
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 79 -2.25
		name groundSlab228
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 76.5 -4.25
		name groundSlab229
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 77.5 -4.25
		name groundSlab230
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 87 -1.75
		name groundSlab231
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 89 -3.75
		name groundSlab233
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 88 -3.75
		name groundSlab234
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 87 -3.75
		name groundSlab235
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 86 -1.75
		name groundSlab236
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 84 -3
		name groundSlab237
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 83 -3
		name groundSlab238
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 82 -3
		name groundSlab239
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 81 -5
		name groundSlab240
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 80 -5
		name groundSlab241
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 2 -1.75
		name groundSlab42
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 0 -3.75
		name groundSlab44
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 1 -3.75
		name groundSlab45
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 2 -3.75
		name groundSlab46
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 3 -1.75
		name groundSlab47
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 5 -3
		name groundSlab48
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 6 -3
		name groundSlab49
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 7 -3
		name groundSlab50
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 8 -5
		name groundSlab51
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 9 -5
		name groundSlab52
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 11.5 -4.25
		name groundSlab55
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 12.5 -4.25
		name groundSlab56
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 10 -2.25
		name groundSlab57
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 12 -0.75
		name groundSlab58
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 13 -0.75
		name groundSlab62
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 14 -0.75
		name groundSlab63
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 15 -0.75
		name groundSlab64
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 16 -0.75
		name groundSlab65
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 17 -0.75
		name groundSlab67
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 17 -0.75
		name groundSlab68
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 19 -2.25
		name groundSlab69
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 16.5 -4.25
		name groundSlab70
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 17.5 -4.25
		name groundSlab71
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 27 -1.75
		name groundSlab72
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 29 -3.75
		name groundSlab74
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 28 -3.75
		name groundSlab75
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 27 -3.75
		name groundSlab76
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 26 -1.75
		name groundSlab77
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 24 -3
		name groundSlab78
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 23 -3
		name groundSlab79
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 22 -3
		name groundSlab80
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 21 -5
		name groundSlab81
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
WorldObject{
	ObjectProperties{
		position 20 -5
		name groundSlab82
		texture slab
	}
	PhysicObjectProperties{
		type static
		shape box
		density 1
		friction 0.3
		angle 0
		velocity 0 0
	}
	WorldObjectProperties{
	}
}
Spawn{
	position 2 -2.5
}
Spawn{
	position 27 -2.5
}
Spawn{
	position 10 -3
}
Spawn{
	position 19 -3
}
Spawn{
	position 32 -2.5
}
Spawn{
	position 57 -2.5
}
Spawn{
	position 40 -3
}
Spawn{
	position 49 -3
}
Spawn{
	position 62 -2.5
}
Spawn{
	position 87 -2.5
}
Spawn{
	position 70 -3
}
Spawn{
	position 79 -3
}
