fireball Assets/Audio/RPG-SFX/spell_02.ogg
magicMissle Assets/Audio/RPG-SFX/spell_01.ogg
arrow Assets/Audio/RPG-SFX/wood_02.ogg
menu Assets/Audio/menu.wav
eqChange Assets/Audio/RPG-SFX/misc_01.ogg
collect Assets/Audio/BonusCube.ogg
jump Assets/Audio/jump.ogg
hit Assets/Audio/RPG-SFX/creature_misc_01.ogg
laserBall Assets/Audio/RPG-SFX/spell_fire_06.ogg