Weapon{
	ObjectProperties{
		position -0.484848 -0.484848
		name bow
		texture bow
	}
	ItemProperties{
		amount 266814656
		isWorldObject true
		textureOnEquip bowEquiped
	}
	WeaponProperties{
		attackDelay 600
		bulletSpeed 1000
		dmg 7
		reloadSpeed 1000
		maxAmmo 1
		ammo 1
		bulletTexture arrow
		bulletDistance 55
		reloading false
		shotSound arrow
	}
}
Weapon{
	ObjectProperties{
		position -0.484848 -0.484848
		name dagger
		texture dagger
	}
	ItemProperties{
		amount 266709088
		isWorldObject true
		textureOnEquip daggerEquiped
	}
	WeaponProperties{
		attackDelay 1000
		bulletSpeed 500
		dmg 100
		reloadSpeed 1000
		maxAmmo 1
		ammo 1
		bulletTexture transparent
		bulletDistance 0.01
		reloading false
		shotSound arrow
	}
}
Weapon{
	ObjectProperties{
		position -0.484848 -0.484848
		name laserRod
		texture laserRod
	}
	ItemProperties{
		amount 266709088
		isWorldObject true
		textureOnEquip laserRodEquiped
	}
	WeaponProperties{
		attackDelay 25
		bulletSpeed 350
		dmg 1
		reloadSpeed 3000
		maxAmmo 50
		ammo 50
		bulletTexture laserBall
		bulletDistance 2
		reloading false
		shotSound laserBall
	}
}
Item{
	ObjectProperties{
		position 0 0
		name nothing
		texture 
	}
	ItemProperties{
		amount 0
		isWorldObject false
		textureOnEquip nothing
	}
}
Weapon{
	ObjectProperties{
		position -0.484848 -0.484848
		name rodBrown
		texture rodBrown
	}
	ItemProperties{
		amount 266709088
		isWorldObject true
		textureOnEquip rodBrownEquiped
	}
	WeaponProperties{
		attackDelay 250
		bulletSpeed 1000
		dmg 2
		reloadSpeed 1000
		maxAmmo 10
		ammo 10
		bulletTexture laser
		bulletDistance 10
		reloading false
		shotSound magicMissle
	}
}
Weapon{
	ObjectProperties{
		position -0.484848 -0.484848
		name staff
		texture staff
	}
	ItemProperties{
		amount 266708992
		isWorldObject true
		textureOnEquip staffRubyEquiped
	}
	WeaponProperties{
		attackDelay 400
		bulletSpeed 1000
		dmg 3
		reloadSpeed 3000
		maxAmmo 20
		ammo 20
		bulletTexture fireball
		bulletDistance 25
		reloading false
		shotSound fireball
	}
}
