Player{
	ObjectProperties{
		position 52.0273 -0.972727
		name player2
		texture humanMale
	}
	PhysicObjectProperties{
		type dynamic
		shape circle
		density 1
		friction 0.1
		angle 0
		velocity 0 0
	}
	EntityProperties{
		maxHP 30
		HP 0
		jumpHeight 300
		movementSpeed 10
		isFacingLeft false
		equiped 0
		EQ{
			rodBrown 10 3733
			bow 1 32833
			nothing 0
			nothing 0
			nothing 0
		}
	}
	PlayerProperties{
		textureBase humanMale
		textureHair aragornHair
		textureBoots bootsMiddleGray
		textureLegs legArmor0
		textureGloves gloveBrown
		textureBody aragornBody
		textureHandRight rodBrownEquiped
		textureCloak cloackBlack
		textureBeard nothing
	}
}
