Weapon{
	ObjectProperties{
		position -0.484848 -0.484848
		name bow
		texture bow
	}
	ItemProperties{
		amount 807405744
		isWorldObject true
		textureOnEquip bowEquiped
	}
	WeaponProperties{
		attackDelay 600
		bulletSpeed 1000
		dmg 7
		reloadSpeed 1200
		maxAmmo 1
		ammo 1
		bulletTexture arrow
		bulletDistance 50
		reloading false
		shotSound arrow
	}
}
Item{
	ObjectProperties{
		position 0 0
		name nothing
		texture 
	}
	ItemProperties{
		amount 0
		isWorldObject false
		textureOnEquip nothing
	}
}
Weapon{
	ObjectProperties{
		position -0.484848 -0.484848
		name rodBrown
		texture rodBrown
	}
	ItemProperties{
		amount 807300176
		isWorldObject true
		textureOnEquip rodBrownEquiped
	}
	WeaponProperties{
		attackDelay 250
		bulletSpeed 1000
		dmg 2
		reloadSpeed 1000
		maxAmmo 10
		ammo 10
		bulletTexture laser
		bulletDistance 15
		reloading false
		shotSound magicMissle
	}
}
Weapon{
	ObjectProperties{
		position -0.484848 -0.484848
		name staff
		texture staff
	}
	ItemProperties{
		amount 807300080
		isWorldObject true
		textureOnEquip staffRubyEquiped
	}
	WeaponProperties{
		attackDelay 350
		bulletSpeed 1000
		dmg 3
		reloadSpeed 3000
		maxAmmo 20
		ammo 20
		bulletTexture fireball
		bulletDistance 30
		reloading false
		shotSound fireball
	}
}
