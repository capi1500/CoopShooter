Weapon{
    ObjectProperties{
        name assultRifle
    }
    ItemProperties{
        ammount 1
        worldObject false
    }
    WeaponProperties{
        attackDelay 250
        bulletSpeed 50
        dmg 2
        reloadSpeed 3000
        maxAmmo 15
        bulletTexture arrow
    }
}
Weapon{
    ObjectProperties{
        name bazooka
    }
    ItemProperties{
        ammount 1
        worldObject false
    }
    WeaponProperties{
        attackDelay 750
        bulletSpeed 15
        dmg 6
        reloadSpeed 2000
        maxAmmo 1
        bulletTexture fireball
    }
}
Weapon{
    ObjectProperties{
        name minigun
    }
    ItemProperties{
        ammount 1
        worldObject false
    }
    WeaponProperties{
        attackDelay 50
        bulletSpeed 50
        dmg 2
        reloadSpeed 3000
        maxAmmo 45
        bulletTexture fireball
    }
}