Player{
	ObjectProperties{
		position 52.1957 -5.95979
		name player2
		texture humanMale
	}
	PhysicObjectProperties{
		type dynamic
		shape circle
		density 1
		friction 0.1
		angle 0
		velocity -20.6338 62.9413
	}
	EntityProperties{
		maxHP 25
		HP 0
		jumpHeight 300
		movementSpeed 10
		isFacingLeft true
		equiped 1
		EQ{
			rodBrown 10 56043
			bow 1 3866
			nothing 0
			nothing 0
			nothing 0
		}
	}
	PlayerProperties{
		textureBase humanMale
		textureHair aragornHair
		textureBoots bootsMiddleGray
		textureLegs legArmor0
		textureGloves gloveBrown
		textureBody aragornBody
		textureHandRight bowEquiped
		textureCloak cloackBlack
		textureBeard nothing
	}
}
