Player{
	ObjectProperties{
		position 47.9727 -0.975305
		name player1
		texture humanMale
	}
	PhysicObjectProperties{
		type dynamic
		shape circle
		density 1
		friction 0.1
		angle 0
		velocity 0 0
	}
	EntityProperties{
		maxHP 25
		HP 5
		jumpHeight 300
		movementSpeed 10
		isFacingLeft true
		equiped 0
		EQ{
			staff 8 32833
			nothing 0
			nothing 0
			nothing 0
			nothing 0
		}
	}
	PlayerProperties{
		textureBase humanMale
		textureHair longWhiteHair
		textureBoots bootsMiddleGray
		textureLegs nothing
		textureGloves nothing
		textureBody gandalfBody
		textureHandRight staffRubyEquiped
		textureCloak cloackGray
		textureBeard nothing
	}
}
