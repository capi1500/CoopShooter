Weapon{
    ObjectProperties{
        name bow
        texture bow
    }
    ItemProperties{
        ammount 1
        worldObject false
        textureOnEquip bowEquiped
    }
    WeaponProperties{
        attackDelay 500
        bulletSpeed 50
        dmg 6
        reloadSpeed 500
        maxAmmo 1
        bulletTexture arrow
        bulletDistance 50
    }
}
Weapon{
    ObjectProperties{
        name rodBrown
        texture rodBrown
    }
    ItemProperties{
        ammount 1
        worldObject false
        textureOnEquip rodBrownEquiped
    }
    WeaponProperties{
        attackDelay 350
        bulletSpeed 50
        dmg 2
        reloadSpeed 3000
        maxAmmo 10
        bulletTexture laser
        bulletDistance 20
    }
}
Weapon{
    ObjectProperties{
        name staff
        texture staff
    }
    ItemProperties{
        ammount 1
        worldObject false
        textureOnEquip staffRubyEquiped
    }
    WeaponProperties{
        attackDelay 300
        bulletSpeed 50
        dmg 2
        reloadSpeed 3000
        maxAmmo 20
        bulletTexture fireball
        bulletDistance 30
    }
}