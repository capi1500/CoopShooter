Weapon{
	ObjectProperties{
		position -1.45455 -1.45455
		name bow
		texture bow
	}
	ItemProperties{
		amount 1
		isWorldObject false
		textureOnEquip bowEquiped
	}
	WeaponProperties{
		attackDelay 500
		bulletSpeed 1000
		dmg 6
		reloadSpeed 500
		maxAmmo 1
		ammo 1
		bulletTexture arrow
		bulletDistance 50
		reloading false
		shotSound arrow
	}
}
Item{
	ObjectProperties{
		position 0 0
		name nothing
		texture }
	}
	ItemProperties{
		amount 1
		isWorldObject false
		textureOnEquip nothing
	}
}
Weapon{
	ObjectProperties{
		position -1.45455 -1.45455
		name rodBrown
		texture rodBrown
	}
	ItemProperties{
		amount -709313616
		isWorldObject true
		textureOnEquip rodBrownEquiped
	}
	WeaponProperties{
		attackDelay 350
		bulletSpeed 1000
		dmg 2
		reloadSpeed 3000
		maxAmmo 10
		ammo 7
		bulletTexture laser
		bulletDistance 20
		reloading false
		shotSound magicMissle
	}
}
Weapon{
	ObjectProperties{
		position -1.45455 -1.45455
		name staff
		texture staff
	}
	ItemProperties{
		amount -709313712
		isWorldObject true
		textureOnEquip staffRubyEquiped
	}
	WeaponProperties{
		attackDelay 300
		bulletSpeed 1000
		dmg 2
		reloadSpeed 3000
		maxAmmo 20
		ammo 20
		bulletTexture fireball
		bulletDistance 30
		reloading false
		shotSound fireball
	}
}
