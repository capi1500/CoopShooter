Player{
	ObjectProperties{
		position 54.214 -0.973754
		name player1
		texture humanMale
	}
	PhysicObjectProperties{
		type dynamic
		shape circle
		density 1
		friction 0.1
		angle 0
		velocity 0 0
	}
	EntityProperties{
		maxHP 30
		HP 16
		jumpHeight 300
		movementSpeed 10
		isFacingLeft false
		equiped 1
		EQ{
			dagger 1 56043
			laserRod 50 3649
			nothing 0
			nothing 0
			nothing 0
		}
	}
	PlayerProperties{
		textureBase humanMale
		textureHair longWhiteHair
		textureBoots bootsMiddleGray
		textureLegs nothing
		textureGloves nothing
		textureBody gandalfBody
		textureHandRight laserRodEquiped
		textureCloak cloackGray
		textureBeard nothing
	}
}
