wall.png box
slab.png slab
ground.png ground
wall.png wall
heal.png healCollect
hpUp.png hpUpCollect
dmgUp.png dmgUpCollect
fasterShots.png fasterShotsCollect
fasterShooting.png fasterShootingCollect
noReload.png noReloadCollect
health.png healthBar
ammo.png ammoBar
battlemage.png mage
archer.png archer
arrow.png arrow
fireball.png fireball