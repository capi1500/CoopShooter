WorldObject{
	ObjectProperties{
	    position 200 5
	    name ground1
	    texture ground
	}
	PhysicObjectProperties{
        shape box
	}
}
WorldObject{
    ObjectProperties{
 	    position 600 5
 	    name ground2
 	    texture ground
	}
	PhysicObjectProperties{
        shape box
	}
}
WorldObject{
    ObjectProperties{
 	    position 1000 5
 	    name ground3
 	    texture ground
	}
	PhysicObjectProperties{
        shape box
	}
}
WorldObject{
	ObjectProperties{
	    position -5 -195
	    name wall1
	    texture wall
	}
	PhysicObjectProperties{
        shape box
	}
}
WorldObject{
	ObjectProperties{
	    position 1205 -195
	    name wall2
	    texture wall
	}
	PhysicObjectProperties{
        shape box
	}
}
WorldObject{
    ObjectProperties{
        position 100 -50
        name box1
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 100 -20
        name box2
        texture box
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 20 -130
        name box3
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 60 -130
        name box4
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 100 -130
        name box5
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 140 -50
        name box6
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 220 -100
        name box7
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position  260 -100
        name box8
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 300 -100
        name box9
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 340 -180
        name box10
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 380 -180
        name box11
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 380 -60
        name box12
        texture box
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 260 -20
        name box13
        texture box
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 480 -150
        name box27
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 520 -150
        name box28
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 420 -70
        name box31
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 500 -10
        name box33
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 540 -80
        name box35
        texture box
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 600 -220
        name box38
        texture box
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 600 -260
        name box37
        texture box
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 540 -10
        name box39
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 580 -10
        name box40
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 620 -10
        name box41
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 660 -10
        name box42
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 660 -80
        name box46
        texture box
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 700 -10
        name box34
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 700 -10
        name box34
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 780 -70
        name box32
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 680 -150
        name box29
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 720 -150
        name box30
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 1100 -50
        name box14
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 1100 -20
        name box15
        texture box
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 1180 -130
        name box16
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 1140 -130
        name box17
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 1100 -130
        name box18
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 1060 -50
        name box19
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 980 -100
        name box20
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 940 -100
        name box21
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 900 -100
        name box22
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 860 -180
        name box23
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 820 -180
        name box24
        texture slab
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 820 -60
        name box25
        texture box
    }
    PhysicObjectProperties{
        shape box
    }
}
WorldObject{
    ObjectProperties{
        position 940 -20
        name box26
        texture box
    }
    PhysicObjectProperties{
        shape box
    }
}