WorldObject{
	ObjectProperties{
	    position 235 465
	    name ground1
	    texture ground
	}
	PhysicObjectProperties{
        shape box
	}
}
WorldObject{
    ObjectProperties{
 	    position 685 465
 	    name ground2
 	    texture ground
	}
	PhysicObjectProperties{
        shape box
	}
}
WorldObject{
    ObjectProperties{
 	    position 1135 465
 	    name ground3
 	    texture ground
	}
	PhysicObjectProperties{
        shape box
	}
}
WorldObject{
	ObjectProperties{
	    position 5 235
	    name wall1
	    texture wall
	}
	PhysicObjectProperties{
        shape box
	}
}
WorldObject{
	ObjectProperties{
	    position 1365 235
	    name wall2
	    texture wall
	}
	PhysicObjectProperties{
        shape box
	}
}