Player{
    ObjectProperties{
        position 1180 -20
        name player2
        texture ballYellow
    }
    PhysicObjectProperties{
        type dynamic
        shape circle
        friction 0.1
        density 1
    }
    EntityProperties{
        maxHP 10
        HP 10
        jumpHeight 300
        movementSpeed 10
        EQ{
            gun 1
        }
    }
}